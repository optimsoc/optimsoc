../system_2x2_cccc/optimsoc_def.vh