`define FLIT32_WIDTH 34
