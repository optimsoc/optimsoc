// Address of the Diagnosis Processor
`define DBG_NOC_ADDR_DP 5'd2


// diagnosis system snapshot packet (from packetizer)
`define DBG_NOC_CLASS_DIAG_SNAPSHOT 3'b110

