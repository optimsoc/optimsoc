../system_2x2_cccc/tb_system_2x2_cccc.sv