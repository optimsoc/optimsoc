../compute_tile/tb_compute_tile.sv