/* Copyright (c) 2013 by the author(s)
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
 * THE SOFTWARE.
 *
 * =============================================================================
 *
 * Cross-Trigger Matrix (CTM)
 *
 * Author(s):
 *   Philipp Wagner <mail@philipp-wagner.com>
 */

`include "dbg_config.vh"

`include "lisnoc_def.vh"
`include "lisnoc16_def.vh"

module ctm(/*AUTOARG*/
   // Outputs
   dbgnoc_out_flit, dbgnoc_out_valid, dbgnoc_in_ready,
   trigger_from_ctm,
   // Inputs
   clk, rst, dbgnoc_out_ready, dbgnoc_in_flit, dbgnoc_in_valid,
   trigger_to_ctm
   );

   // parameters for the Debug NoC interface
   parameter DBG_NOC_DATA_WIDTH = `FLIT16_CONTENT_WIDTH;
   parameter DBG_NOC_FLIT_TYPE_WIDTH = `FLIT16_TYPE_WIDTH;
   localparam DBG_NOC_FLIT_WIDTH = DBG_NOC_DATA_WIDTH + DBG_NOC_FLIT_TYPE_WIDTH;
   parameter DBG_NOC_PH_DEST_WIDTH = `FLIT16_DEST_WIDTH;
   parameter DBG_NOC_PH_CLASS_WIDTH = `PACKET16_CLASS_WIDTH;
   localparam DBG_NOC_PH_ID_WIDTH = DBG_NOC_DATA_WIDTH - DBG_NOC_PH_DEST_WIDTH - DBG_NOC_PH_CLASS_WIDTH;
   parameter DBG_NOC_VCHANNELS = 'hx;

   // number of debug module
   parameter DEBUG_MODULE_COUNT = 'hx;

   // module description
   localparam MODULE_TYPE_CTM = 8'h01;
   localparam MODULE_VERSION_CTM = 8'h00;

   // number of configuration registers required to hold all cross-trigger
   // configuration entries (one bit per input trigger)
   // ceil(DEBUG_MODULE_COUNT/16) with integers
   localparam TRIGGER_CONF_REGISTERS = 1 + ((DEBUG_MODULE_COUNT - 1) / 16);

   localparam CONF_MEM_SIZE = 1 + TRIGGER_CONF_REGISTERS;

   input clk;
   input rst;

   // Debug NoC interface (IN = NoC -> CTM; OUT = CTM -> NoC)
   output [DBG_NOC_FLIT_WIDTH-1:0] dbgnoc_out_flit;
   output [DBG_NOC_VCHANNELS-1:0] dbgnoc_out_valid;
   input [DBG_NOC_VCHANNELS-1:0] dbgnoc_out_ready;
   input [DBG_NOC_FLIT_WIDTH-1:0] dbgnoc_in_flit;
   input [DBG_NOC_VCHANNELS-1:0] dbgnoc_in_valid;
   output [DBG_NOC_VCHANNELS-1:0] dbgnoc_in_ready;

   // trigger interface
   output [DEBUG_MODULE_COUNT-1:0] trigger_from_ctm;
   input [DEBUG_MODULE_COUNT-1:0] trigger_to_ctm;

   wire [DEBUG_MODULE_COUNT-1:0] conf_triggers_enabled;

   // Right now all trigger outputs get the same trigger signal.
   // For eventual forward compatibility we leave the multiple trigger outputs
   // in place.
   wire trigger_from_ctm_single;
   assign trigger_from_ctm = {DEBUG_MODULE_COUNT{trigger_from_ctm_single}};

   // configuration memory
   wire [CONF_MEM_SIZE*16-1:0] conf_mem_flat_in;
   reg [CONF_MEM_SIZE-1:0] conf_mem_flat_in_valid;
   wire [CONF_MEM_SIZE*16-1:0] conf_mem_flat_out;

   // un-flatten conf_mem_in to conf_mem_flat_in
   reg [15:0] conf_mem_in [CONF_MEM_SIZE-1:0];
   genvar i;
   generate
      for (i = 0; i < CONF_MEM_SIZE; i = i + 1) begin : gen_conf_mem_in
         assign conf_mem_flat_in[((i+1)*16)-1:i*16] = conf_mem_in[i];
      end
   endgenerate

   // un-flatten conf_mem_flat_out to conf_mem_out
   wire [15:0] conf_mem_out [CONF_MEM_SIZE-1:0];
   generate
      for (i = 0; i < CONF_MEM_SIZE; i = i + 1) begin : gen_conf_mem_out
         assign conf_mem_out[i] = conf_mem_flat_out[((i+1)*16)-1:i*16];
      end
   endgenerate

   /* dbgnoc_conf_if AUTO_TEMPLATE(
      .dbgnoc_out_rts(),
      .conf_mem_flat_in_ack(),
      .\(.*\)(\1), // suppress explict port widths
    ); */
   dbgnoc_conf_if
      #(.MEM_SIZE(CONF_MEM_SIZE),
        .MEM_INIT_ZERO(0))
      u_dbgnoc_conf_if(/*AUTOINST*/
                       // Outputs
                       .dbgnoc_out_flit (dbgnoc_out_flit),       // Templated
                       .dbgnoc_out_valid(dbgnoc_out_valid),      // Templated
                       .dbgnoc_in_ready (dbgnoc_in_ready),       // Templated
                       .dbgnoc_out_rts  (),                      // Templated
                       .conf_mem_flat_out(conf_mem_flat_out),    // Templated
                       .conf_mem_flat_in_ack(),                  // Templated
                       // Inputs
                       .clk             (clk),                   // Templated
                       .rst             (rst),                   // Templated
                       .dbgnoc_out_ready(dbgnoc_out_ready),      // Templated
                       .dbgnoc_in_flit  (dbgnoc_in_flit),        // Templated
                       .dbgnoc_in_valid (dbgnoc_in_valid),       // Templated
                       .conf_mem_flat_in(conf_mem_flat_in),      // Templated
                       .conf_mem_flat_in_valid(conf_mem_flat_in_valid)); // Templated

   // configuration register initialization
   always @ (posedge clk) begin
      if (rst) begin
         // initialize configuration registers
         conf_mem_in[0] = {MODULE_TYPE_CTM, MODULE_VERSION_CTM};
         // all other registers are set to 0 in the generate block below
         conf_mem_flat_in_valid <= {CONF_MEM_SIZE{1'b1}};
      end else begin
         conf_mem_flat_in_valid <= 0;
      end
   end

   generate
      for (i = 1; i < 1 + TRIGGER_CONF_REGISTERS; i = i + 1) begin
         always @ (posedge clk) begin
            if (rst) begin
               conf_mem_in[i] <= 0; // disable all cross-triggers by default
            end
         end
      end
   endgenerate

   // build a conf_triggers_enabled signal out of the individual configuration
   // registers
   genvar j;
   generate
      for (i = 1; i < 1 + TRIGGER_CONF_REGISTERS; i = i + 1) begin
         for (j = 0; j < 16; j = j + 1) begin
            if ((i-1)*16 + j < DEBUG_MODULE_COUNT) begin
               assign conf_triggers_enabled[(i-1)*16 + j] = conf_mem_out[i][j];
            end
         end
      end
   endgenerate

   // triggering
   assign trigger_from_ctm_single =| (conf_triggers_enabled & trigger_to_ctm);

endmodule
