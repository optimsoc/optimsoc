../compute_tile/optimsoc_def.vh